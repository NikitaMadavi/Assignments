magic
tech sky130A
timestamp 1726418409
<< error_p >>
rect 432 50 506 68
rect 432 23 450 50
rect 488 23 506 50
rect 432 5 506 23
<< nwell >>
rect -301 584 449 586
rect -465 495 554 584
rect -464 195 554 495
rect -301 193 449 195
<< nmos >>
rect -390 15 -375 150
rect -30 14 -1 60
rect 180 14 211 60
rect 390 14 421 60
<< pmos >>
rect -390 254 -375 435
rect -30 389 -1 435
rect 180 389 211 435
rect 390 389 421 435
<< ndiff >>
rect -435 120 -390 150
rect -435 45 -427 120
rect -402 45 -390 120
rect -435 15 -390 45
rect -375 120 -330 150
rect -375 45 -367 120
rect -342 45 -330 120
rect -375 15 -330 45
rect -135 14 -30 60
rect -1 14 180 60
rect 211 14 390 60
rect 421 50 509 60
rect 421 23 450 50
rect 488 23 509 50
rect 421 14 509 23
<< pdiff >>
rect -435 375 -390 435
rect -435 315 -426 375
rect -400 315 -390 375
rect -435 254 -390 315
rect -375 375 -330 435
rect -120 389 -30 435
rect -1 389 180 435
rect 211 389 390 435
rect 421 389 508 435
rect -375 315 -364 375
rect -338 315 -330 375
rect -375 254 -330 315
<< ndiffc >>
rect -427 45 -402 120
rect -367 45 -342 120
<< pdiffc >>
rect -426 315 -400 375
rect -364 315 -338 375
<< psubdiff >>
rect -436 -61 -331 -44
rect -436 -90 -405 -61
rect -359 -90 -331 -61
rect -436 -105 -331 -90
<< nsubdiff >>
rect -427 540 -338 560
rect -427 509 -407 540
rect -360 509 -338 540
rect -427 486 -338 509
rect 450 23 488 50
<< psubdiffcont >>
rect -405 -90 -359 -61
<< nsubdiffcont >>
rect -407 509 -360 540
<< poly >>
rect -390 435 -375 464
rect -30 435 -1 464
rect 180 435 211 464
rect 390 435 421 465
rect -390 150 -375 254
rect -30 60 -1 389
rect 180 60 211 389
rect 390 60 421 389
rect -390 -15 -375 15
rect -30 -15 -1 14
rect 180 -15 211 14
rect 390 -14 421 14
<< locali >>
rect -421 540 -346 549
rect -421 509 -407 540
rect -360 509 -346 540
rect -421 499 -346 509
rect -431 375 -396 390
rect -431 315 -426 375
rect -400 315 -396 375
rect -431 300 -396 315
rect -369 375 -334 390
rect -369 315 -364 375
rect -338 315 -334 375
rect -369 300 -334 315
rect -431 120 -398 135
rect -431 45 -427 120
rect -402 45 -398 120
rect -431 30 -398 45
rect -371 120 -338 135
rect -371 45 -367 120
rect -342 45 -338 120
rect -371 30 -338 45
rect -420 -61 -345 -54
rect -420 -90 -405 -61
rect -359 -90 -345 -61
rect -420 -97 -345 -90
<< viali >>
rect -397 516 -371 533
rect -397 -86 -366 -66
<< metal1 >>
rect -555 533 375 539
rect -555 516 -397 533
rect -371 516 375 533
rect -555 511 375 516
rect -555 510 -211 511
rect -526 -66 479 -61
rect -526 -86 -397 -66
rect -366 -86 479 -66
rect -526 -91 479 -86
<< labels >>
rlabel metal1 -282 527 -282 527 1 VDD
<< end >>
