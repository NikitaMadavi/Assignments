magic
tech sky130A
timestamp 1726399087
<< locali >>
rect 615 395 665 405
rect 615 390 625 395
rect -100 370 0 390
rect 320 370 625 390
rect 615 365 625 370
rect 655 365 665 395
rect 615 355 665 365
rect 1775 395 1825 405
rect 1775 365 1785 395
rect 1815 390 1825 395
rect 1815 370 1990 390
rect 1815 365 1825 370
rect 1775 355 1825 365
rect -100 130 0 150
rect 460 130 685 150
rect 1665 130 1990 150
rect 2450 130 2700 150
rect 3680 130 3880 150
rect 685 50 705 130
rect 520 30 705 50
rect -100 10 0 30
rect 285 -200 305 0
rect 405 -200 445 -190
rect 285 -220 415 -200
rect 435 -220 445 -200
rect 405 -230 445 -220
rect 520 -440 540 30
rect 615 0 665 10
rect 615 -30 625 0
rect 655 -5 665 0
rect 1715 0 1760 10
rect 1715 -5 1725 0
rect 655 -25 1725 -5
rect 1750 -25 1760 0
rect 655 -30 665 -25
rect 615 -40 665 -30
rect 1715 -35 1760 -25
rect 645 -200 685 -190
rect 1775 -195 1825 -185
rect 1775 -200 1785 -195
rect 645 -220 655 -200
rect 675 -220 960 -200
rect 1280 -220 1785 -200
rect 645 -230 685 -220
rect 1775 -225 1785 -220
rect 1815 -225 1825 -195
rect 1775 -235 1825 -225
rect 1900 -440 1920 130
rect 1990 0 2035 10
rect 1990 -25 2000 0
rect 2025 -25 2035 0
rect 1990 -35 2035 -25
rect 2275 -180 2295 0
rect 1970 -195 2020 -185
rect 1970 -225 1980 -195
rect 2010 -200 2020 -195
rect 2260 -190 2310 -180
rect 2010 -220 2185 -200
rect 2010 -225 2020 -220
rect 1970 -235 2020 -225
rect 520 -460 960 -440
rect 1420 -460 1920 -440
rect 2165 -560 2185 -220
rect 2260 -220 2270 -190
rect 2300 -220 2310 -190
rect 2260 -230 2310 -220
rect 2770 -440 2790 130
rect 2820 -190 2870 -180
rect 2820 -220 2830 -190
rect 2860 -200 2870 -190
rect 2860 -220 2990 -200
rect 2820 -230 2870 -220
rect 3560 -265 3610 -255
rect 3560 -295 3570 -265
rect 3600 -295 3610 -265
rect 3560 -305 3610 -295
rect 3735 -265 3785 -255
rect 3735 -295 3745 -265
rect 3775 -295 3785 -265
rect 3735 -305 3785 -295
rect 3830 -440 3850 130
rect 2770 -460 2990 -440
rect 3450 -460 3850 -440
rect 2165 -580 2990 -560
rect 1245 -620 1265 -590
rect 2260 -615 2310 -605
rect 2260 -620 2270 -615
rect 1245 -640 2270 -620
rect 2260 -645 2270 -640
rect 2300 -645 2310 -615
rect 2260 -655 2310 -645
<< viali >>
rect 625 365 655 395
rect 1785 365 1815 395
rect 415 -220 435 -200
rect 625 -30 655 0
rect 1725 -25 1750 0
rect 655 -220 675 -200
rect 1785 -225 1815 -195
rect 2000 -25 2025 0
rect 1980 -225 2010 -195
rect 2270 -220 2300 -190
rect 2830 -220 2860 -190
rect 3570 -295 3600 -265
rect 3745 -295 3775 -265
rect 2270 -645 2300 -615
<< metal1 >>
rect 615 395 665 405
rect 615 365 625 395
rect 655 365 665 395
rect 615 355 665 365
rect 1775 395 1825 405
rect 1775 365 1785 395
rect 1815 365 1825 395
rect 1775 355 1825 365
rect -100 205 0 320
rect 145 205 165 320
rect 460 205 685 315
rect 1665 205 1990 315
rect 2135 205 2155 320
rect 2450 205 2700 315
rect 3680 220 3770 240
rect -100 60 0 95
rect 200 60 220 95
rect 460 65 685 95
rect 1665 65 1990 95
rect 2190 60 2210 95
rect 2450 65 2705 95
rect 615 0 665 10
rect 615 -30 625 0
rect 655 -30 665 0
rect 615 -40 665 -30
rect 1715 0 1760 10
rect 1715 -25 1725 0
rect 1750 -5 1760 0
rect 1990 0 2035 10
rect 1990 -5 2000 0
rect 1750 -25 2000 -5
rect 2025 -25 2035 0
rect 1715 -35 1760 -25
rect 1990 -35 2035 -25
rect 405 -200 445 -190
rect 645 -200 685 -190
rect 405 -220 415 -200
rect 435 -220 655 -200
rect 675 -220 685 -200
rect 405 -230 445 -220
rect 645 -230 685 -220
rect 1775 -195 1825 -185
rect 1775 -225 1785 -195
rect 1815 -225 1825 -195
rect 1775 -235 1825 -225
rect 1970 -195 2020 -185
rect 1970 -225 1980 -195
rect 2010 -225 2020 -195
rect 1970 -235 2020 -225
rect 2260 -190 2310 -180
rect 2260 -220 2270 -190
rect 2300 -220 2310 -190
rect 2260 -230 2310 -220
rect 2820 -190 2870 -180
rect 2820 -220 2830 -190
rect 2860 -220 2870 -190
rect 2820 -230 2870 -220
rect 3560 -265 3610 -255
rect 3560 -270 3570 -265
rect 1105 -385 1125 -270
rect 1420 -385 2990 -270
rect 3135 -385 3155 -270
rect 3450 -295 3570 -270
rect 3600 -295 3610 -265
rect 3560 -305 3610 -295
rect 3660 -495 3680 65
rect 3750 -255 3770 220
rect 3735 -265 3785 -255
rect 3735 -295 3745 -265
rect 3775 -295 3785 -265
rect 3735 -305 3785 -295
rect 1160 -530 1180 -495
rect 1420 -530 2990 -495
rect 3190 -530 3210 -495
rect 3450 -530 3680 -495
rect 2260 -615 2310 -605
rect 2260 -645 2270 -615
rect 2300 -645 2310 -615
rect 2260 -655 2310 -645
<< via1 >>
rect 625 365 655 395
rect 1785 365 1815 395
rect 625 -30 655 0
rect 1785 -225 1815 -195
rect 1980 -225 2010 -195
rect 2270 -220 2300 -190
rect 2830 -220 2860 -190
rect 3570 -295 3600 -265
rect 3745 -295 3775 -265
rect 2270 -645 2300 -615
<< metal2 >>
rect 615 395 665 405
rect 615 365 625 395
rect 655 365 665 395
rect 615 355 665 365
rect 1775 395 1825 405
rect 1775 365 1785 395
rect 1815 365 1825 395
rect 1775 355 1825 365
rect 630 10 650 355
rect 615 0 665 10
rect 615 -30 625 0
rect 655 -30 665 0
rect 615 -40 665 -30
rect 1790 -185 1810 355
rect 1775 -195 1825 -185
rect 1775 -225 1785 -195
rect 1815 -200 1825 -195
rect 1970 -195 2020 -185
rect 1970 -200 1980 -195
rect 1815 -220 1980 -200
rect 1815 -225 1825 -220
rect 1775 -235 1825 -225
rect 1970 -225 1980 -220
rect 2010 -225 2020 -195
rect 1970 -235 2020 -225
rect 2260 -190 2310 -180
rect 2260 -220 2270 -190
rect 2300 -195 2310 -190
rect 2820 -190 2870 -180
rect 2820 -195 2830 -190
rect 2300 -215 2830 -195
rect 2300 -220 2310 -215
rect 2260 -230 2310 -220
rect 2820 -220 2830 -215
rect 2860 -220 2870 -190
rect 2820 -230 2870 -220
rect 2275 -605 2295 -230
rect 3560 -265 3610 -255
rect 3560 -295 3570 -265
rect 3600 -270 3610 -265
rect 3735 -265 3785 -255
rect 3735 -270 3745 -265
rect 3600 -295 3745 -270
rect 3775 -295 3785 -265
rect 3560 -305 3610 -295
rect 3735 -305 3785 -295
rect 2260 -615 2310 -605
rect 2260 -645 2270 -615
rect 2300 -645 2310 -615
rect 2260 -655 2310 -645
use inverter  inverter_0
timestamp 1726254829
transform 1 0 995 0 1 55
box -310 -10 180 300
use inverter  inverter_1
timestamp 1726254829
transform 1 0 1485 0 1 55
box -310 -10 180 300
use inverter  inverter_2
timestamp 1726254829
transform 1 0 3010 0 1 55
box -310 -10 180 300
use inverter  inverter_3
timestamp 1726254829
transform 1 0 3500 0 1 55
box -310 -10 180 300
use tg1  tg1_0
timestamp 1726394591
transform 1 0 1250 0 1 -550
box -290 -40 170 355
use tg1  tg1_1
timestamp 1726394591
transform 1 0 2280 0 1 40
box -290 -40 170 355
use tg  tg_0
timestamp 1726394604
transform 1 0 290 0 1 40
box -290 -40 170 355
use tg  tg_1
timestamp 1726394604
transform 1 0 3280 0 1 -550
box -290 -40 170 355
<< labels >>
flabel locali -100 140 -100 140 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali 3880 140 3880 140 0 FreeSans 400 0 0 0 Q
port 2 nsew
flabel locali -100 20 -100 20 0 FreeSans 400 0 0 0 clk
port 3 nsew
flabel locali -100 380 -100 380 0 FreeSans 400 0 0 0 clk_bar
port 4 nsew
flabel metal1 -100 260 -100 260 0 FreeSans 400 0 0 0 vdd
port 5 nsew
flabel metal1 -100 75 -100 75 0 FreeSans 400 0 0 0 vss
port 7 nsew
<< end >>
