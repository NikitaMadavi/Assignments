VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dff2
  CLASS BLOCK ;
  FOREIGN dff2 ;
  ORIGIN 1.000 6.550 ;
  SIZE 39.800 BY 10.600 ;
  PIN D
    ANTENNADIFFAREA 2.182500 ;
    PORT
      LAYER li1 ;
        RECT 1.650 2.050 2.800 3.200 ;
        RECT 2.200 1.500 2.400 2.050 ;
        RECT -1.000 1.300 2.400 1.500 ;
        RECT 2.200 0.950 2.400 1.300 ;
        RECT 2.200 0.600 2.800 0.950 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA 4.365000 ;
    PORT
      LAYER li1 ;
        RECT 35.250 2.000 36.350 3.150 ;
        RECT 35.650 1.500 35.850 2.000 ;
        RECT 35.650 1.300 38.800 1.500 ;
        RECT 35.650 1.000 35.850 1.300 ;
        RECT 35.250 0.650 35.850 1.000 ;
        RECT 33.050 -3.850 34.200 -2.700 ;
        RECT 33.450 -4.400 33.650 -3.850 ;
        RECT 38.300 -4.400 38.500 1.300 ;
        RECT 33.450 -4.600 38.500 -4.400 ;
        RECT 33.450 -4.950 33.650 -4.600 ;
        RECT 33.050 -5.300 33.650 -4.950 ;
    END
  END Q
  PIN clk
    ANTENNAGATEAREA 0.540000 ;
    PORT
      LAYER li1 ;
        RECT 17.750 3.900 18.250 4.050 ;
        RECT 22.650 3.900 23.100 3.950 ;
        RECT 17.750 3.700 23.100 3.900 ;
        RECT 17.750 3.550 18.250 3.700 ;
        RECT 22.650 3.550 23.100 3.700 ;
        RECT 2.750 0.300 3.200 0.400 ;
        RECT -1.000 0.100 3.200 0.300 ;
        RECT 2.750 0.000 3.200 0.100 ;
        RECT 2.850 -2.000 3.050 0.000 ;
        RECT 4.050 -2.000 4.450 -1.900 ;
        RECT 2.850 -2.200 4.450 -2.000 ;
        RECT 4.050 -2.300 4.450 -2.200 ;
        RECT 6.450 -2.000 6.850 -1.900 ;
        RECT 12.350 -2.000 12.800 -1.950 ;
        RECT 17.750 -2.000 18.250 -1.850 ;
        RECT 6.450 -2.200 18.250 -2.000 ;
        RECT 6.450 -2.300 6.850 -2.200 ;
        RECT 12.350 -2.350 12.800 -2.200 ;
        RECT 17.750 -2.350 18.250 -2.200 ;
        RECT 19.700 -2.000 20.200 -1.850 ;
        RECT 19.700 -2.200 21.850 -2.000 ;
        RECT 19.700 -2.350 20.200 -2.200 ;
        RECT 21.650 -5.600 21.850 -2.200 ;
        RECT 32.650 -5.600 33.100 -5.500 ;
        RECT 21.650 -5.800 33.100 -5.600 ;
        RECT 32.650 -5.900 33.100 -5.800 ;
      LAYER met1 ;
        RECT 17.750 3.550 18.250 4.050 ;
        RECT 4.050 -2.000 4.450 -1.900 ;
        RECT 6.450 -2.000 6.850 -1.900 ;
        RECT 4.050 -2.200 6.850 -2.000 ;
        RECT 4.050 -2.300 4.450 -2.200 ;
        RECT 6.450 -2.300 6.850 -2.200 ;
        RECT 17.750 -2.350 18.250 -1.850 ;
        RECT 19.700 -2.350 20.200 -1.850 ;
      LAYER met2 ;
        RECT 17.750 3.550 18.250 4.050 ;
        RECT 17.900 -1.850 18.100 3.550 ;
        RECT 17.750 -2.000 18.250 -1.850 ;
        RECT 19.700 -2.000 20.200 -1.850 ;
        RECT 17.750 -2.200 20.200 -2.000 ;
        RECT 17.750 -2.350 18.250 -2.200 ;
        RECT 19.700 -2.350 20.200 -2.200 ;
    END
  END clk
  PIN clk_bar
    ANTENNAGATEAREA 0.540000 ;
    PORT
      LAYER li1 ;
        RECT 2.750 3.900 3.200 3.950 ;
        RECT 6.150 3.900 6.650 4.050 ;
        RECT -1.000 3.700 6.650 3.900 ;
        RECT 2.750 3.550 3.200 3.700 ;
        RECT 6.150 3.550 6.650 3.700 ;
        RECT 22.650 0.300 23.100 0.400 ;
        RECT 19.900 0.100 23.100 0.300 ;
        RECT 6.150 -0.050 6.650 0.100 ;
        RECT 17.150 -0.050 17.600 0.100 ;
        RECT 6.150 -0.250 17.600 -0.050 ;
        RECT 6.150 -0.400 6.650 -0.250 ;
        RECT 17.150 -0.350 17.600 -0.250 ;
        RECT 19.900 -0.350 20.350 0.100 ;
        RECT 22.650 0.000 23.100 0.100 ;
        RECT 22.750 -1.800 22.950 0.000 ;
        RECT 22.600 -2.300 23.100 -1.800 ;
        RECT 28.200 -2.000 28.700 -1.800 ;
        RECT 32.650 -2.000 33.100 -1.950 ;
        RECT 28.200 -2.200 33.100 -2.000 ;
        RECT 28.200 -2.300 28.700 -2.200 ;
        RECT 32.650 -2.350 33.100 -2.200 ;
        RECT 12.350 -5.600 12.800 -5.500 ;
        RECT 9.600 -5.800 12.800 -5.600 ;
        RECT 12.350 -5.900 12.800 -5.800 ;
        RECT 12.450 -6.200 12.650 -5.900 ;
        RECT 22.600 -6.200 23.100 -6.050 ;
        RECT 12.450 -6.400 23.100 -6.200 ;
        RECT 22.600 -6.550 23.100 -6.400 ;
      LAYER met1 ;
        RECT 6.150 3.550 6.650 4.050 ;
        RECT 6.150 -0.400 6.650 0.100 ;
        RECT 17.150 -0.050 17.600 0.100 ;
        RECT 19.900 -0.050 20.350 0.100 ;
        RECT 17.150 -0.250 20.350 -0.050 ;
        RECT 17.150 -0.350 17.600 -0.250 ;
        RECT 19.900 -0.350 20.350 -0.250 ;
        RECT 22.600 -2.300 23.100 -1.800 ;
        RECT 28.200 -2.300 28.700 -1.800 ;
        RECT 22.600 -6.550 23.100 -6.050 ;
      LAYER met2 ;
        RECT 6.150 3.550 6.650 4.050 ;
        RECT 6.300 0.100 6.500 3.550 ;
        RECT 6.150 -0.400 6.650 0.100 ;
        RECT 22.600 -1.950 23.100 -1.800 ;
        RECT 28.200 -1.950 28.700 -1.800 ;
        RECT 22.600 -2.150 28.700 -1.950 ;
        RECT 22.600 -2.300 23.100 -2.150 ;
        RECT 28.200 -2.300 28.700 -2.150 ;
        RECT 22.750 -6.050 22.950 -2.300 ;
        RECT 22.600 -6.550 23.100 -6.050 ;
    END
  END clk_bar
  PIN vdd
    ANTENNADIFFAREA 21.869999 ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.750 4.600 3.500 ;
        RECT 6.850 1.700 16.650 3.550 ;
        RECT 19.900 1.750 24.500 3.500 ;
        RECT 27.000 1.700 36.800 3.550 ;
        RECT 9.600 -4.150 14.200 -2.400 ;
        RECT 29.900 -4.150 34.500 -2.400 ;
      LAYER li1 ;
        RECT 0.300 2.050 1.450 3.200 ;
        RECT 7.350 2.000 9.850 3.150 ;
        RECT 12.250 2.000 14.750 3.150 ;
        RECT 20.200 2.050 21.350 3.200 ;
        RECT 27.500 2.000 30.000 3.150 ;
        RECT 32.400 2.000 34.900 3.150 ;
        RECT 9.900 -3.850 11.050 -2.700 ;
        RECT 30.200 -3.850 31.350 -2.700 ;
        RECT 35.600 -3.050 36.100 -2.550 ;
        RECT 37.350 -3.050 37.850 -2.550 ;
      LAYER met1 ;
        RECT -1.000 3.150 4.600 3.200 ;
        RECT 19.900 3.150 24.500 3.200 ;
        RECT -1.000 2.400 36.800 3.150 ;
        RECT -1.000 2.200 37.700 2.400 ;
        RECT -1.000 2.050 36.800 2.200 ;
        RECT 6.850 2.000 16.650 2.050 ;
        RECT 27.000 2.000 36.800 2.050 ;
        RECT 37.500 -2.550 37.700 2.200 ;
        RECT 35.600 -2.700 36.100 -2.550 ;
        RECT 9.600 -2.950 36.100 -2.700 ;
        RECT 9.600 -3.850 34.500 -2.950 ;
        RECT 35.600 -3.050 36.100 -2.950 ;
        RECT 37.350 -3.050 37.850 -2.550 ;
      LAYER met2 ;
        RECT 35.600 -2.700 36.100 -2.550 ;
        RECT 37.350 -2.700 37.850 -2.550 ;
        RECT 35.600 -2.950 37.850 -2.700 ;
        RECT 35.600 -3.050 36.100 -2.950 ;
        RECT 37.350 -3.050 37.850 -2.950 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER li1 ;
        RECT 1.400 0.600 2.000 0.950 ;
        RECT 8.450 0.650 9.850 1.000 ;
        RECT 13.350 0.650 14.750 1.000 ;
        RECT 21.300 0.600 21.900 0.950 ;
        RECT 28.600 0.650 30.000 1.000 ;
        RECT 33.500 0.650 34.900 1.000 ;
        RECT 11.000 -5.300 11.600 -4.950 ;
        RECT 31.300 -5.300 31.900 -4.950 ;
      LAYER met1 ;
        RECT 6.850 0.950 16.650 1.000 ;
        RECT 27.000 0.950 36.800 1.000 ;
        RECT -1.000 0.650 36.800 0.950 ;
        RECT -1.000 0.600 4.600 0.650 ;
        RECT 19.900 0.600 24.500 0.650 ;
        RECT 36.600 -4.950 36.800 0.650 ;
        RECT 9.600 -5.300 36.800 -4.950 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 3.150 2.050 4.300 3.200 ;
        RECT 3.550 1.500 3.750 2.050 ;
        RECT 10.200 2.000 11.300 3.150 ;
        RECT 15.100 2.000 16.200 3.150 ;
        RECT 21.550 2.050 22.700 3.200 ;
        RECT 23.050 2.050 24.200 3.200 ;
        RECT 9.550 1.500 9.950 1.600 ;
        RECT 3.550 1.300 9.950 1.500 ;
        RECT 3.550 0.950 3.750 1.300 ;
        RECT 3.150 0.600 3.750 0.950 ;
        RECT 6.850 0.500 7.050 1.300 ;
        RECT 9.550 1.200 9.950 1.300 ;
        RECT 10.600 1.500 10.800 2.000 ;
        RECT 14.450 1.500 14.850 1.600 ;
        RECT 10.600 1.300 14.850 1.500 ;
        RECT 10.600 1.000 10.800 1.300 ;
        RECT 14.450 1.200 14.850 1.300 ;
        RECT 15.500 1.500 15.700 2.000 ;
        RECT 22.100 1.500 22.300 2.050 ;
        RECT 15.500 1.300 22.300 1.500 ;
        RECT 15.500 1.000 15.700 1.300 ;
        RECT 10.200 0.650 10.800 1.000 ;
        RECT 15.100 0.650 15.700 1.000 ;
        RECT 5.200 0.300 7.050 0.500 ;
        RECT 5.200 -4.400 5.400 0.300 ;
        RECT 11.250 -3.850 12.400 -2.700 ;
        RECT 12.750 -3.850 13.900 -2.700 ;
        RECT 11.800 -4.400 12.000 -3.850 ;
        RECT 5.200 -4.600 12.000 -4.400 ;
        RECT 11.800 -4.950 12.000 -4.600 ;
        RECT 13.150 -4.400 13.350 -3.850 ;
        RECT 19.000 -4.400 19.200 1.300 ;
        RECT 22.100 0.950 22.300 1.300 ;
        RECT 23.450 1.500 23.650 2.050 ;
        RECT 30.350 2.000 31.450 3.150 ;
        RECT 29.700 1.500 30.100 1.600 ;
        RECT 23.450 1.300 30.100 1.500 ;
        RECT 23.450 0.950 23.650 1.300 ;
        RECT 22.100 0.600 22.700 0.950 ;
        RECT 23.050 0.600 23.650 0.950 ;
        RECT 13.150 -4.600 19.200 -4.400 ;
        RECT 27.700 -4.400 27.900 1.300 ;
        RECT 29.700 1.200 30.100 1.300 ;
        RECT 30.750 1.500 30.950 2.000 ;
        RECT 34.600 1.500 35.000 1.600 ;
        RECT 30.750 1.300 35.000 1.500 ;
        RECT 30.750 1.000 30.950 1.300 ;
        RECT 34.600 1.200 35.000 1.300 ;
        RECT 30.350 0.650 30.950 1.000 ;
        RECT 31.550 -3.850 32.700 -2.700 ;
        RECT 32.100 -4.400 32.300 -3.850 ;
        RECT 27.700 -4.600 32.300 -4.400 ;
        RECT 13.150 -4.950 13.350 -4.600 ;
        RECT 11.800 -5.300 12.400 -4.950 ;
        RECT 12.750 -5.300 13.350 -4.950 ;
        RECT 32.100 -4.950 32.300 -4.600 ;
        RECT 32.100 -5.300 32.700 -4.950 ;
  END
END dff2
END LIBRARY

