MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.980 0.250 ;
  SIZE 1.980 BY 3.000 ;
  PIN A
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT -0.550 0.620 0.000 0.870 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 0.528000 ;
    PORT
      LAYER li1 ;
        RECT 0.230 0.820 0.400 2.460 ;
        RECT 0.230 0.650 0.860 0.820 ;
        RECT 0.230 0.000 0.400 0.650 ;
    END
  END Y
  PIN vdd
    ANTENNADIFFAREA 1.072000 ;
    PORT
      LAYER nwell ;
        RECT -0.980 0.940 0.630 2.640 ;
      LAYER li1 ;
        RECT -0.600 2.580 -0.200 2.720 ;
        RECT -0.750 1.120 -0.080 2.580 ;
      LAYER met1 ;
        RECT -0.800 2.500 0.950 2.750 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 0.315000 ;
    PORT
      LAYER li1 ;
        RECT -0.650 -0.150 -0.080 0.420 ;
      LAYER met1 ;
        RECT -0.750 -0.250 1.000 0.050 ;
    END
  END vss
END INVX1
END LIBRARY

