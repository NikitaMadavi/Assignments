* Nikita Suresh Madavi
* 23M1160
* Negative edge D flipflop

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Subcircuit definition of inverter
.subckt inverter A Y vdd vss
XMP1 Y A vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.34 ad=.402 as=.402 pd=3.28 ps=3.28
XMN1 Y A vss vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.45 ad=0.135 as=0.135 pd=1.5 ps=1.5
.ends inverter

* Subcircuit definition of transmission gate
.subckt tg D Q clk clk_bar vdd vss
XMP2 D clk_bar Q vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.34 ad=.402 as=.402 pd=3.28 ps=3.28
XMN2 D clk Q vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.45 ad=0.135 as=0.135 pd=1.5 ps=1.5
.ends tg

* Subcircuit definition of transmission gate
.subckt tg1 D Q clk clk_bar vdd vss
XMP3 D clk Q vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.34 ad=.402 as=.402 pd=3.28 ps=3.28
XMN4 D clk_bar Q vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.45 ad=0.135 as=0.135 pd=1.5 ps=1.5
.ends tg1

* D flipflop defination
.subckt dff D Q clk clk_bar vdd vss
Xtg1 D q1 clk clk_bar vdd vss tg

Xinv1 q1 qn vdd vss inverter
Xinv2 qn q2 vdd vss inverter
Xtg2 q2 qn clk_bar clk vdd vss tg1

Xtg3 q2 q3 clk_bar clk vdd vss tg1

Xinv3 q3 q4 vdd vss inverter
Xinv4 q4 Q vdd vss inverter
Xtg4 Q q4 clk clk_bar vdd vss tg
.ends dff

Xd1 D Q clk clk_bar vdd vss dff



