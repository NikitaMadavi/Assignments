magic
tech sky130A
timestamp 1725804771
<< nwell >>
rect -98 94 63 264
<< nmos >>
rect 0 0 15 42
<< pmos >>
rect 0 112 15 246
<< ndiff >>
rect -30 30 0 42
rect -30 10 -25 30
rect -8 10 0 30
rect -30 0 0 10
rect 15 30 45 42
rect 15 10 23 30
rect 40 10 45 30
rect 15 0 45 10
<< pdiff >>
rect -30 217 0 246
rect -30 142 -25 217
rect -8 142 0 217
rect -30 112 0 142
rect 15 217 45 246
rect 15 142 23 217
rect 40 142 45 217
rect 15 112 45 142
<< ndiffc >>
rect -25 10 -8 30
rect 23 10 40 30
<< pdiffc >>
rect -25 142 -8 217
rect 23 142 40 217
<< psubdiff >>
rect -75 30 -30 42
rect -75 10 -60 30
rect -43 10 -30 30
rect -75 0 -30 10
<< nsubdiff >>
rect -80 217 -30 246
rect -80 142 -70 217
rect -53 142 -30 217
rect -80 112 -30 142
<< psubdiffcont >>
rect -60 10 -43 30
<< nsubdiffcont >>
rect -70 142 -53 217
<< poly >>
rect 0 246 15 259
rect 0 89 15 112
rect -36 84 15 89
rect -36 67 -25 84
rect -8 67 15 84
rect -36 60 15 67
rect 0 42 15 60
rect 0 -13 15 0
<< polycont >>
rect -25 67 -8 84
<< locali >>
rect -75 255 -60 258
rect -20 255 -8 258
rect -75 217 -8 255
rect -75 142 -70 217
rect -53 142 -25 217
rect -75 112 -8 142
rect 23 217 40 246
rect -55 84 0 87
rect -55 67 -25 84
rect -8 67 0 84
rect -55 62 0 67
rect 23 82 40 142
rect 23 65 86 82
rect -65 30 -8 42
rect -65 10 -60 30
rect -43 10 -25 30
rect -65 2 -8 10
rect -65 -15 -45 2
rect -25 -15 -8 2
rect 23 30 40 65
rect 23 0 40 10
<< viali >>
rect -60 255 -20 272
rect -45 -15 -25 2
<< metal1 >>
rect -80 272 95 275
rect -80 255 -60 272
rect -20 255 95 272
rect -80 250 95 255
rect -75 2 100 5
rect -75 -15 -45 2
rect -25 -15 100 2
rect -75 -25 100 -15
<< labels >>
rlabel locali -55 75 -55 75 7 A
port 1 w
rlabel locali 86 75 86 75 3 Y
port 2 e
rlabel metal1 95 265 95 265 3 vdd
port 3 e
rlabel metal1 100 -10 100 -10 3 vss
port 4 e
<< end >>
